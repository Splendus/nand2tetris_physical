/**
 * Not gate:
 * out = not in
 */

`default_nettype none
module Not(
	input in,
	output out
);
    
    Nand(out,in,in); 

endmodule
